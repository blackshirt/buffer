module buffer

import math 

const (
	max_buffer_size = math.max_u16
)
